module FP16MAC(
  input  [7:0] io_a,
  input  [7:0] io_b,
  input  [7:0] io_c,
  output [7:0] io_out
);
  wire [15:0] _io_out_T = io_a * io_b; // @[PE_INT8.scala 11:19]
  wire [15:0] _GEN_0 = {{8'd0}, io_c}; // @[PE_INT8.scala 11:27]
  wire [15:0] _io_out_T_2 = _io_out_T + _GEN_0; // @[PE_INT8.scala 11:27]
  assign io_out = _io_out_T_2[7:0]; // @[PE_INT8.scala 11:10]
endmodule
module FP16PE(
  input        clock,
  input        reset,
  input  [7:0] io_vecA_0,
  input  [7:0] io_vecA_1,
  input  [7:0] io_vecA_2,
  input  [7:0] io_vecA_3,
  input  [7:0] io_vecA_4,
  input  [7:0] io_vecA_5,
  input  [7:0] io_vecA_6,
  input  [7:0] io_vecA_7,
  input  [7:0] io_vecA_8,
  input  [7:0] io_vecA_9,
  input  [7:0] io_vecA_10,
  input  [7:0] io_vecA_11,
  input  [7:0] io_vecA_12,
  input  [7:0] io_vecA_13,
  input  [7:0] io_vecA_14,
  input  [7:0] io_vecA_15,
  input  [7:0] io_vecB_0,
  input  [7:0] io_vecB_1,
  input  [7:0] io_vecB_2,
  input  [7:0] io_vecB_3,
  input  [7:0] io_vecB_4,
  input  [7:0] io_vecB_5,
  input  [7:0] io_vecB_6,
  input  [7:0] io_vecB_7,
  input  [7:0] io_vecB_8,
  input  [7:0] io_vecB_9,
  input  [7:0] io_vecB_10,
  input  [7:0] io_vecB_11,
  input  [7:0] io_vecB_12,
  input  [7:0] io_vecB_13,
  input  [7:0] io_vecB_14,
  input  [7:0] io_vecB_15,
  output [7:0] io_resultMAC
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] macs_0_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_0_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_0_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_0_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_1_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_1_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_1_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_1_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_2_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_2_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_2_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_2_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_3_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_3_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_3_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_3_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_4_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_4_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_4_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_4_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_5_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_5_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_5_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_5_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_6_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_6_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_6_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_6_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_7_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_7_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_7_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_7_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_8_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_8_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_8_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_8_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_9_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_9_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_9_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_9_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_10_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_10_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_10_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_10_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_11_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_11_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_11_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_11_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_12_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_12_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_12_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_12_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_13_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_13_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_13_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_13_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_14_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_14_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_14_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_14_io_out; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_15_io_a; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_15_io_b; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_15_io_c; // @[PE_INT8.scala 22:33]
  wire [7:0] macs_15_io_out; // @[PE_INT8.scala 22:33]
  reg [7:0] accumulator_0; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_1; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_2; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_3; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_4; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_5; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_6; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_7; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_8; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_9; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_10; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_11; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_12; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_13; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_14; // @[PE_INT8.scala 25:28]
  reg [7:0] accumulator_15; // @[PE_INT8.scala 25:28]
  FP16MAC macs_0 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_0_io_a),
    .io_b(macs_0_io_b),
    .io_c(macs_0_io_c),
    .io_out(macs_0_io_out)
  );
  FP16MAC macs_1 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_1_io_a),
    .io_b(macs_1_io_b),
    .io_c(macs_1_io_c),
    .io_out(macs_1_io_out)
  );
  FP16MAC macs_2 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_2_io_a),
    .io_b(macs_2_io_b),
    .io_c(macs_2_io_c),
    .io_out(macs_2_io_out)
  );
  FP16MAC macs_3 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_3_io_a),
    .io_b(macs_3_io_b),
    .io_c(macs_3_io_c),
    .io_out(macs_3_io_out)
  );
  FP16MAC macs_4 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_4_io_a),
    .io_b(macs_4_io_b),
    .io_c(macs_4_io_c),
    .io_out(macs_4_io_out)
  );
  FP16MAC macs_5 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_5_io_a),
    .io_b(macs_5_io_b),
    .io_c(macs_5_io_c),
    .io_out(macs_5_io_out)
  );
  FP16MAC macs_6 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_6_io_a),
    .io_b(macs_6_io_b),
    .io_c(macs_6_io_c),
    .io_out(macs_6_io_out)
  );
  FP16MAC macs_7 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_7_io_a),
    .io_b(macs_7_io_b),
    .io_c(macs_7_io_c),
    .io_out(macs_7_io_out)
  );
  FP16MAC macs_8 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_8_io_a),
    .io_b(macs_8_io_b),
    .io_c(macs_8_io_c),
    .io_out(macs_8_io_out)
  );
  FP16MAC macs_9 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_9_io_a),
    .io_b(macs_9_io_b),
    .io_c(macs_9_io_c),
    .io_out(macs_9_io_out)
  );
  FP16MAC macs_10 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_10_io_a),
    .io_b(macs_10_io_b),
    .io_c(macs_10_io_c),
    .io_out(macs_10_io_out)
  );
  FP16MAC macs_11 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_11_io_a),
    .io_b(macs_11_io_b),
    .io_c(macs_11_io_c),
    .io_out(macs_11_io_out)
  );
  FP16MAC macs_12 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_12_io_a),
    .io_b(macs_12_io_b),
    .io_c(macs_12_io_c),
    .io_out(macs_12_io_out)
  );
  FP16MAC macs_13 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_13_io_a),
    .io_b(macs_13_io_b),
    .io_c(macs_13_io_c),
    .io_out(macs_13_io_out)
  );
  FP16MAC macs_14 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_14_io_a),
    .io_b(macs_14_io_b),
    .io_c(macs_14_io_c),
    .io_out(macs_14_io_out)
  );
  FP16MAC macs_15 ( // @[PE_INT8.scala 22:33]
    .io_a(macs_15_io_a),
    .io_b(macs_15_io_b),
    .io_c(macs_15_io_c),
    .io_out(macs_15_io_out)
  );
  assign io_resultMAC = accumulator_15; // @[PE_INT8.scala 37:16]
  assign macs_0_io_a = io_vecA_0; // @[PE_INT8.scala 27:18]
  assign macs_0_io_b = io_vecB_0; // @[PE_INT8.scala 28:18]
  assign macs_0_io_c = 8'h0; // @[PE_INT8.scala 29:18]
  assign macs_1_io_a = io_vecA_1; // @[PE_INT8.scala 32:22]
  assign macs_1_io_b = io_vecB_1; // @[PE_INT8.scala 33:22]
  assign macs_1_io_c = accumulator_0; // @[PE_INT8.scala 34:22]
  assign macs_2_io_a = io_vecA_2; // @[PE_INT8.scala 32:22]
  assign macs_2_io_b = io_vecB_2; // @[PE_INT8.scala 33:22]
  assign macs_2_io_c = accumulator_1; // @[PE_INT8.scala 34:22]
  assign macs_3_io_a = io_vecA_3; // @[PE_INT8.scala 32:22]
  assign macs_3_io_b = io_vecB_3; // @[PE_INT8.scala 33:22]
  assign macs_3_io_c = accumulator_2; // @[PE_INT8.scala 34:22]
  assign macs_4_io_a = io_vecA_4; // @[PE_INT8.scala 32:22]
  assign macs_4_io_b = io_vecB_4; // @[PE_INT8.scala 33:22]
  assign macs_4_io_c = accumulator_3; // @[PE_INT8.scala 34:22]
  assign macs_5_io_a = io_vecA_5; // @[PE_INT8.scala 32:22]
  assign macs_5_io_b = io_vecB_5; // @[PE_INT8.scala 33:22]
  assign macs_5_io_c = accumulator_4; // @[PE_INT8.scala 34:22]
  assign macs_6_io_a = io_vecA_6; // @[PE_INT8.scala 32:22]
  assign macs_6_io_b = io_vecB_6; // @[PE_INT8.scala 33:22]
  assign macs_6_io_c = accumulator_5; // @[PE_INT8.scala 34:22]
  assign macs_7_io_a = io_vecA_7; // @[PE_INT8.scala 32:22]
  assign macs_7_io_b = io_vecB_7; // @[PE_INT8.scala 33:22]
  assign macs_7_io_c = accumulator_6; // @[PE_INT8.scala 34:22]
  assign macs_8_io_a = io_vecA_8; // @[PE_INT8.scala 32:22]
  assign macs_8_io_b = io_vecB_8; // @[PE_INT8.scala 33:22]
  assign macs_8_io_c = accumulator_7; // @[PE_INT8.scala 34:22]
  assign macs_9_io_a = io_vecA_9; // @[PE_INT8.scala 32:22]
  assign macs_9_io_b = io_vecB_9; // @[PE_INT8.scala 33:22]
  assign macs_9_io_c = accumulator_8; // @[PE_INT8.scala 34:22]
  assign macs_10_io_a = io_vecA_10; // @[PE_INT8.scala 32:22]
  assign macs_10_io_b = io_vecB_10; // @[PE_INT8.scala 33:22]
  assign macs_10_io_c = accumulator_9; // @[PE_INT8.scala 34:22]
  assign macs_11_io_a = io_vecA_11; // @[PE_INT8.scala 32:22]
  assign macs_11_io_b = io_vecB_11; // @[PE_INT8.scala 33:22]
  assign macs_11_io_c = accumulator_10; // @[PE_INT8.scala 34:22]
  assign macs_12_io_a = io_vecA_12; // @[PE_INT8.scala 32:22]
  assign macs_12_io_b = io_vecB_12; // @[PE_INT8.scala 33:22]
  assign macs_12_io_c = accumulator_11; // @[PE_INT8.scala 34:22]
  assign macs_13_io_a = io_vecA_13; // @[PE_INT8.scala 32:22]
  assign macs_13_io_b = io_vecB_13; // @[PE_INT8.scala 33:22]
  assign macs_13_io_c = accumulator_12; // @[PE_INT8.scala 34:22]
  assign macs_14_io_a = io_vecA_14; // @[PE_INT8.scala 32:22]
  assign macs_14_io_b = io_vecB_14; // @[PE_INT8.scala 33:22]
  assign macs_14_io_c = accumulator_13; // @[PE_INT8.scala 34:22]
  assign macs_15_io_a = io_vecA_15; // @[PE_INT8.scala 32:22]
  assign macs_15_io_b = io_vecB_15; // @[PE_INT8.scala 33:22]
  assign macs_15_io_c = accumulator_14; // @[PE_INT8.scala 34:22]
  always @(posedge clock) begin
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_0 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_0 <= macs_0_io_out; // @[PE_INT8.scala 30:20]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_1 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_1 <= macs_1_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_2 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_2 <= macs_2_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_3 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_3 <= macs_3_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_4 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_4 <= macs_4_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_5 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_5 <= macs_5_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_6 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_6 <= macs_6_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_7 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_7 <= macs_7_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_8 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_8 <= macs_8_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_9 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_9 <= macs_9_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_10 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_10 <= macs_10_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_11 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_11 <= macs_11_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_12 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_12 <= macs_12_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_13 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_13 <= macs_13_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_14 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_14 <= macs_14_io_out; // @[PE_INT8.scala 35:24]
    end
    if (reset) begin // @[PE_INT8.scala 25:28]
      accumulator_15 <= 8'h0; // @[PE_INT8.scala 25:28]
    end else begin
      accumulator_15 <= macs_15_io_out; // @[PE_INT8.scala 35:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  accumulator_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  accumulator_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  accumulator_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  accumulator_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  accumulator_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  accumulator_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  accumulator_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  accumulator_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  accumulator_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  accumulator_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  accumulator_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  accumulator_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  accumulator_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  accumulator_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  accumulator_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  accumulator_15 = _RAND_15[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
